library ieee;
use ieee.std_logic_1164.all;

entity OutputBufferControl_tb is
end OutputBufferControl_tb;

architecture behavioral of OutputBufferControl_tb is

    -- Componente a testar
    component OutputBufferControl is
        port (
            reset   : in  std_logic;
            clk     : in  std_logic;
            Load    : in  std_logic;
            ACK     : in  std_logic;
            Wreg    : out std_logic;
            OBfree  : out std_logic;
            Dval    : out std_logic
        );
    end component;

    -- Constantes de tempo
    constant clk_period      : time := 10 ns;
    constant half_clk_period : time := clk_period / 2;

    -- Sinais de estímulo e observação
    signal clk_tb     : std_logic;
    signal reset_tb   : std_logic;
    signal Load_tb    : std_logic;
    signal ACK_tb     : std_logic;
    signal Wreg_tb    : std_logic;
    signal OBfree_tb  : std_logic;
    signal Dval_tb    : std_logic;

begin

    -- Instância do DUT
    UUT: OutputBufferControl
        port map (
            reset   => reset_tb,
            clk     => clk_tb,
            Load    => Load_tb,
            ACK     => ACK_tb,
            Wreg    => Wreg_tb,
            OBfree  => OBfree_tb,
            Dval    => Dval_tb
        );

    -- Clock generator
    clk_gen: process
    begin
        while true loop
            clk_tb <= '0';
            wait for half_clk_period;
            clk_tb <= '1';
            wait for half_clk_period;
        end loop;
    end process;

    -- Estímulos para percorrer todos os estados
    stimulus: process
    begin
        -- RESET para garantir estado inicial
        reset_tb <= '1';
		  ACK_tb   <= '0';
		  Load_tb  <= '0';
        wait for clk_period;
        reset_tb <= '0';
        wait for clk_period;

        -- Estado Idle → Load → WaitAck → Clear → Idle

        -- S1: Ativar Load para passar de Idle para Load
        Load_tb <= '1';
        wait for clk_period;

        -- S2: Desativar Load (transição para WaitAck ocorre mesmo assim)
        Load_tb <= '0';
        wait for clk_period;

        -- S3: Manter em WaitAck, ACK = 0 (ficar no mesmo estado)
        wait for clk_period;

        -- S4: Enviar ACK → transição para Clear
        ACK_tb <= '1';
        wait for clk_period;

        -- S5: Desativar ACK → Clear → Idle
        ACK_tb <= '0';
        wait for clk_period;

        -- Repetição opcional para robustez (nova carga)
        Load_tb <= '1';
        wait for clk_period;
        Load_tb <= '0';
        wait for clk_period;

        ACK_tb <= '1';
        wait for clk_period;
        ACK_tb <= '0';
        wait for clk_period;

        -- Fim da simulação
        wait for clk_period * 3;
    end process;

end behavioral;
