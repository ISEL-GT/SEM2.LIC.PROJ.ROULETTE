LIBRARY ieee: 
USE ieee.std_logic_1164.all;


-- This is the top-level entity responsible for running the actual program
entity roulette is

	port (


	);
		
end roulette;
