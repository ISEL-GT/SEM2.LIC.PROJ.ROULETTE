    Mac OS X            	   2   �      �                                      ATTR       �   �   <                  �   <  com.apple.quarantine q/0083;67b35cdd;Safari;1A25B813-2BE4-413F-B92F-CFAED58B9025 