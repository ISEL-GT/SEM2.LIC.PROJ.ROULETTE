component ficheiro2 is
port (	
	CLK : in std_logic;
	RESET : in std_logic;
	SET : in std_logic;
	D : in std_logic;
	EN : in std_logic;
	Q : out std_logic);
end component;