LIBRARY ieee;
USE ieee.std_logic_1164.all;


-- This is the top-level entity responsible for running the actual program
entity key_decode_rtb is

	port (
		Kack 	: 	in std_logic;
		lines: 	in std_logic_vector(3 downto 0);
		CLK	:	in std_logic;
		Reset :	in std_logic;

		columns : 	out std_logic_vector(3 downto 0);
		Kout 	: 	out std_logic_vector(3 downto 0);
		Kval 	: 	out std_logic
	);

end key_decode_rtb;

architecture structural of key_decode_rtb is

	component key_decode is
		port (
			Kack 	: 	in std_logic;
			lines: 	in std_logic_vector(3 downto 0);
			CLK	:	in std_logic;
			Reset:	in std_logic;

			columns : 	out std_logic_vector(3 downto 0);
			Kout 	: 	out std_logic_vector(3 downto 0);
			Kval 	: 	out std_logic
		);
	end component;

begin

	instance_key_decode: key_decode
		port map (
			Kack 	=> Kack,
			lines => lines,
			CLK 	=> CLK,
			Reset 	=> Reset,

			columns 	=> columns,
			Kout 	=> Kout,
			Kval 	=> Kval
		);

end structural;