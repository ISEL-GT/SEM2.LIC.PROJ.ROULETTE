library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity counter_tb is
end counter_tb;

architecture behavioral of counter_tb is

    component counter is
        port (
            CE                  : in std_logic;
            CLK                 : in std_logic;
            reset               : in std_logic;
            parallel_load_flag  : in std_logic;
            parallel_load_value : in std_logic_vector(1 downto 0);
            count               : out std_logic_vector(1 downto 0)
        );
    end component;
    
    constant clk_period       : TIME := 10 ns;
    constant half_clk_period  : TIME := clk_period / 2;
    
    signal CE_tb                  : std_logic;
    signal CLK_tb                 : std_logic;
    signal reset_tb               : std_logic;
    signal parallel_load_flag_tb  : std_logic;
    signal parallel_load_value_tb : std_logic_vector(1 downto 0);
    signal count_tb               : std_logic_vector(1 downto 0);
    
begin
    
    UUT: counter
        port map (
            CE                  => CE_tb,
            CLK                 => CLK_tb,
            reset               => reset_tb,
            parallel_load_flag  => parallel_load_flag_tb,
            parallel_load_value => parallel_load_value_tb,
            count               => count_tb
        );
    
    -- Clock Generation
    clk_gen: process
    begin
        while true loop
            CLK_tb <= '0';
            wait for half_clk_period;
            CLK_tb <= '1';
            wait for half_clk_period;
        end loop;
    end process;
    
    -- Stimulus Process
    stimulus: process
    begin
        -- Reset the counter and enable counting
        reset_tb 	<= '1';
		  CE_tb 		<= '1';
		  -- Signal to use on mux that selects the parallel load
		  parallel_load_flag_tb <= '0';
		  -- Value that will be input in the register if the selector is 1
        parallel_load_value_tb <= "01";
        wait for clk_period;
		
        reset_tb 	<= '0';
		  wait for clk_period*8;
		 
              
        parallel_load_flag_tb <= '1';
        wait for clk_period*2;
        
		  -- Stop the increment of the counter by changing the mux signal
        parallel_load_flag_tb <= '1';
		  parallel_load_value_tb <= "10";
		  
        wait for clk_period;
        wait for clk_period;
		  
		  -- Change it to the default form of the counter, increment +1
		  parallel_load_flag_tb <= '0';
		  parallel_load_value_tb <= "01";
			
		  wait for clk_period*8;
        
        -- Disable counting
        CE_tb <= '0';
        wait for clk_period;
        
        wait;
    end process;
    
end behavioral;
