    Mac OS X            	   2   �                                           ATTR         �   L                  �     com.apple.lastuseddate#PS       �   <  com.apple.quarantine +�g    ��;    q/0083;67124be0;Safari;D6C13142-F010-42A0-901E-0CB4D817745D 