library ieee;
use ieee.std_logic_1164.all;

entity roulette_tb is
end roulette_tb;

architecture behavioral of roulette_tb is

    component roulette is 
        port (
            	Liness: 	in std_logic_vector(3 downto 0);
					CLK   :	in std_logic;
					Reset :	in std_logic;		
					
					LCD_RS	: 	out std_logic;
					LCD_EN	: 	out std_logic;			
					LCD_DATA	: 	out std_logic_vector(7 downto 4);
					
					Colss 	: 	out std_logic_vector(3 downto 0);
					Kout  	: 	out std_logic_vector(3 downto 0);
					Kval		: 	out std_logic 
        );
    end component;
    
    constant clk_period       : TIME := 20 ns;
    constant half_clk_period  : TIME := clk_period / 2;
    
	 
    signal lines_tb     : std_logic_vector(3 downto 0);
    signal clk_tb       : std_logic;
    signal reset_tb     : std_logic;
	 
	 signal LCD_RS_tb		: std_logic;
	 signal LCD_EN_tb		: std_logic;
	 signal LCD_DATA_tb	: std_logic_vector(7 downto 4);
	 
	 
	 
    signal columns_tb   : std_logic_vector(3 downto 0);
    signal K_tb         : std_logic_vector(3 downto 0);
    signal Kval_tb      : std_logic;

begin
    
    UUT : roulette 
        port map (            
            Liness	=> lines_tb, 
            CLK   	=> clk_tb, 
            Reset		=> reset_tb, 
				
				LCD_RS	=> LCD_RS_tb,
				LCD_EN	=> LCD_EN_tb,
				LCD_DATA => LCD_DATA_tb,
				
				
            Colss  	=> columns_tb, 
            Kval   	=> Kval_tb, 
            Kout   	=> K_tb
        );
    
    clk_gen: process
    begin
        clk_tb <= '0';
        wait for half_clk_period;
        clk_tb <= '1';
        wait for half_clk_period;
    end process;
    
    stimulus: process
    begin
        reset_tb <= '1';
		  lines_tb <= "1111";		  
        wait for clk_period;
		  		  
        lines_tb <= "1111";  -- not Kpress
        reset_tb <= '0';
        wait for clk_period * 10;

        -- Test of first line
        lines_tb <= "0111";
        wait for clk_period * 10;
        
        
        lines_tb <= "1111";  -- not Kpress
        wait for clk_period * 10;
        
        -- Test of second line
        lines_tb <= "1011";
        wait for clk_period * 10;
        
        lines_tb <= "1111";  -- not Kpress
        wait for clk_period * 10;
        

        -- Test of third line
        lines_tb <= "1101";
        wait for clk_period * 10;
		  
        lines_tb <= "1111";  -- not Kpress
        wait for clk_period * 10;

        -- Test of fourth line
        lines_tb <= "1110";
        wait for clk_period * 10;
        
    
        lines_tb <= "1111";  -- not Kpress
        wait for clk_period * 10;
        

        wait;
    end process;
    
end behavioral;
